netcdf test_atomic_types {
variables:
  byte v8;
  short v16;
  int v32;
  float vf; 
  double vd; 
  char vc;
data:
  v8 = -128;
  v16 = -32768;
  v32 = 2147483647;
  vf = 3.1415926535897932384626433832795;
  vd = 3.141592653589793238462643383279502884197169399375105820974944592;
  vc = '@';
}
