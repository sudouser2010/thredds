netcdf test_atomic_array {
dimensions:
  d1 = 1;
  d2 = 2;
  d3 = 3;
  d4 = 4;
  d5 = 5;
variables:
  short v16(d4);
  double vd(d2);
  char vc(d2);

data:
 v16 = 1, 2, 3, 4 ;
 vd = 17.9, 1024.8 ;
 vc = '@', '&' ;
}
