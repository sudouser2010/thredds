netcdf test_fill {
variables:
  byte v8;
  short v16;
  int v32;
	v32:_FillValue=17;
data:
  v8 = 127;
  v16 = 32700;
  v32 = 111000;
}
