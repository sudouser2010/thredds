netcdf test_atomic_types {
variables:
  byte v8;
  ubyte vu8;
  short v16;
  ushort vu16;
  int v32;
  uint vu32;
  int64 v64;
  uint64 vu64;
  float vf; 
  double vd; 
  char vc;
  string vs;
data:
  v8 = -128;
  vu8 = 255;
  v16 = -32768;
  vu16 = 65535;
  v32 = 2147483647;
  vu32 = 4294967295;
  v64 = 9223372036854775807;
  vu64 = 18446744073709551615;
  vf = 3.1415926535897932384626433832795;
  vd = 3.141592653589793238462643383279502884197169399375105820974944592;
  vc = '@';
  vs = "hello\tworld";
}
